LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE my_data_types IS
    TYPE array2D32 IS ARRAY (NATURAL RANGE <>) OF STD_LOGIC_VECTOR(31 downto 0);
END PACKAGE my_data_types;
